package types;
parameter NUM_ALUs=3;
parameter NUM_Threads=4;
endpackage
