package types;
parameter NUM_ALUs=2;
parameter NUM_Threads=4;
endpackage
