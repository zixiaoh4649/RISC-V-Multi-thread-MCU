package types;
parameter NUM_ALUs=4;
parameter NUM_Threads=4;
endpackage
